module findhit (
    input  logic iV,
    input  logic [3:0]  itag1,
    input  logic [3:0]  itag2,
    output logic  oHit
);
always_comb begin
    
end 

endmodule
