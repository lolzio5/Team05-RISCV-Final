module AluOpForwarderE(
  input  logic [1:0]  iForwardAluOp1,
  input  logic [1:0]  iForwardAluOp2,
  input  logic [31:0] iResultDataW,
  input  logic [31:0] iAluResultOutM,
  input  logic [31:0] iRegData1E,
  input  logic [31:0] iRegData2E,

  output logic [31:0] oAluOp1,
  output logic [31:0] oAluOp2,
);


endmodule